library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

package sprites is

 type slika30x30 is array (0 to 29) of unsigned(29 downto 0);
 constant zoga: slika30x30 := ( 
"000000000000000000000000000000",
"000000000011111111111000000000",
"000000001111111111111110000000",
"000000011111111111111111000000",
"000001111111111111111111110000",
"000011111111111111111111111000",
"000011111111111111111111111000",
"000111111111111111111111111100",
"001111111111111111111111111110",
"001111111111111111111111111110",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"011111111111111111111111111111",
"001111111111111111111111111110",
"001111111111111111111111111110",
"000111111111111111111111111100",
"000011111111111111111111111000",
"000011111111111111111111111000",
"000001111111111111111111110000",
"000000011111111111111111000000",
"000000001111111111111110000000",
"000000000011111111111000000000" ); 

 type slika8x8 is array (0 to 7) of unsigned(7 downto 0); 
 constant lab: slika8x8:= (
 "01011100",
 "01000100",
 "00010000",
 "00111100",
 "00000001",
 "10000001",
 "10001001",
 "00111100" );
 
  type tarca20x79 is array (0 to 19) of unsigned(78 downto 0); 
 constant tarca: tarca20x79:= (
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111");
 
  type srce10x16 is array (0 to 9) of unsigned(15 downto 0); 
 constant srce: srce10x16:= (
 "0011100000111100",
 "0111111011111111",
 "1111111111111111",
 "1111111111111111",
 "0111111111111100",
 "0011111111111000",
 "0001111111110000",
 "0000111111100000",
 "0000011111000000",
 "0000001110000000");
 
end sprites;

